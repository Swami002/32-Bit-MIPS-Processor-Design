module tb_mips32;
    reg clk, reset;
    MIPS32 uut(clk, reset);

    initial begin
        $dumpfile("dump.vcd");
        $dumpvars(0, tb_mips32);
    end

    initial begin
        clk = 0;
        forever #5 clk = ~clk;
    end

    initial begin
        reset = 1; #10;
        reset = 0;

        #200;
        $finish;
    end
endmodule
